module mkreq();

endmodules