module ibse();

endmodule