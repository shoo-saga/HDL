module arb(input ack0,ack1,ack2,ack3, output req0,req1,req2,req3);


endmodule