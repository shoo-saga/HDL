module mkwe();

endmodule